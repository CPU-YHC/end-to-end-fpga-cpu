`timescale 1ns / 1ps

module IO_Controller(

    );
endmodule
